module main

interface Object {
	fn hit(r Ray) []Vec
}

// []Vec