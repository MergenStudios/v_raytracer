module main

// for working with colors
// struct Color